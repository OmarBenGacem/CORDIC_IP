module stage_2();

input clk;
input clk_en;
input rst;
input x_one;
input x_two;
input start
output reg done;
output reg result;
output reg valid;



endmodule