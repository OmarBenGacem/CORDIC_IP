module reg_one_to_two ();

endmodule