module stage_2();



endmodule