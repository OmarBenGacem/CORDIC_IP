module stage_4();

input clk;
input rst;
input clk_en;
input val_1;
input val_2;
input current_val;


endmodule