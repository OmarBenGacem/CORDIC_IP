module reg_two_to_three();


endmodule