module cordic_stage();



endmodule